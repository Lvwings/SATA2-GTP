`define ALIGN        	32'h 7B4A4ABC
`define CONT         	32'h 9999AA7C
`define DMAT         	32'h 3636B57C
`define EOF          	32'h D5D5B57C
`define HOLD         	32'h D5D5AA7C
`define HOLDA        	32'h 9595AA7C
`define PMACK        	32'h 9595957C
`define PMNAK        	32'h F5F5957C
`define PMREQ_P      	32'h 1717B57C
`define PMREQ_S      	32'h 7575957C
`define R_ERR        	32'h 5656B57C
`define R_IP         	32'h 5555B57C
`define R_OK         	32'h 3535B57C
`define R_RDY        	32'h 4A4A957C
`define SOF          	32'h 3737B57C
`define SYNC         	32'h B5B5957C
`define WTRM         	32'h 5858B57C
`define X_RDY        	32'h 5757B57C

`define D102			32'h 4A4A4A4A